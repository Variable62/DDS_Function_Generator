module DDS_Top (
    input       wire    Ext_CLK;
    input       wire    Ext_RESETn;
    
);
    
endmodule
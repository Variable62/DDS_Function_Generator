module DDS_Top (

);
end module